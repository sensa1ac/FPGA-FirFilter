module FirFilter 
	#(
		parameter WIDTH = 16, // ширина шины данных
		parameter SIZE =115  // кол-во коэфф-тов КИХ-фильтра (=> и кол-во регистров под отсчёты сигнала x (delay) )
	)
(
	input clk,
	input [WIDTH-1:0] x, // значение текущего отсчёта входного сигнала
	output [WIDTH-1:0]y//output [WIDTH-1:0] y // значение текущего отсчёта выходного сигнала
);
	//wire [WIDTH-1:0] y;
	//assign ty = y[15:0];


	reg [WIDTH-1:0] delay [0:SIZE-1]; // регистры сдвига под отсчеты сигнала x
	wire [WIDTH:0] coef [0:SIZE-1];
	wire [WIDTH-1:0] sum [0:SIZE-1];
	wire [WIDTH-1:0] multres [0:SIZE-1];
	 
		
	// Реализация сдвигового регистра размером SIZE под отсчёты входного сигнала х  
		// На каждый (кроме 1ого) регистр значеине отсчёта идёт с предыдущего
	genvar i;
	generate for(i = SIZE-1; i>0; i=i-1)
	begin: shift
			always @(posedge clk)
			begin	
				delay[i] = delay[i-1];
			end
	end endgenerate	
		// На первый регистр значение отсчёта идёт со входа
	always @(posedge clk)
	begin
		delay[0] = x;
	end
	
	// Реализация SIZE блоков умножителей чисел с фиксированной точкой (рез-т в прямом коде)
	genvar k;
	generate for(k = SIZE-1; k>=0; k=k-1)
	begin: multiply
	multFixPoint #(.Q (WIDTH-2),.N (WIDTH)) // N бит - всё число, Q бит - под дробн. часть
	(
		.mul1(delay[k]), 
		.temp_mul2(coef[k]), 
		.result(multres[k])
	);
	end endgenerate
	
	
	// Итоговое суммирование всех умножений 
	assign sum[0] = multres[0]+multres[1];
	genvar j;
	generate
	for (j = SIZE-1; j>1; j=j-1)
	begin: gensum
		assign sum[j-1] = sum[j-2]+multres[j];
	end
	endgenerate
	
	//*
	/// ???
		d2p d2p1_fir
		(
			.x(y1), 
			.y(y)
		);
	/// ???
	//*/
	
	wire [15:0]y1;
	assign y1 = sum[SIZE-2]; // -2 , т.к. без multres[j], ведь это не итоговая сумма, а только выход из последнего сумматора


// Коэффициенты КИХ-фильтра	часть процесса прямой код   8k 51 ФНЧ 80Дб
/*
assign coef[0] = 17'b10000000000000010;
assign coef[1] = 17'b10000000000001101;
assign coef[2] = 17'b10000000000100011;
assign coef[3] = 17'b10000000001000011;
assign coef[4] = 17'b10000000001100000;
assign coef[5] = 17'b10000000001100110;
assign coef[6] = 17'b10000000001000100;
assign coef[7] = 17'b00000000000000001;
assign coef[8] = 17'b00000000001001001;
assign coef[9] = 17'b00000000001100111;
assign coef[10] = 17'b00000000000111100;
assign coef[11] = 17'b10000000000101000;
assign coef[12] = 17'b10000000010000110;
assign coef[13] = 17'b10000000010010000;
assign coef[14] = 17'b10000000000100111;
assign coef[15] = 17'b00000000010000010;
assign coef[16] = 17'b00000000011110110;
assign coef[17] = 17'b00000000011000000;
assign coef[18] = 17'b10000000000101111;
assign coef[19] = 17'b10000000101010111;
assign coef[20] = 17'b10000000111010110;
assign coef[21] = 17'b10000000011100110;
assign coef[22] = 17'b00000000110011101;
assign coef[23] = 17'b00000010011110111;
assign coef[24] = 17'b00000011111010100;
assign coef[25] = 17'b00000100011110100;
assign coef[26] = 17'b00000011111010100;
assign coef[27] = 17'b00000010011110111;
assign coef[28] = 17'b00000000110011101;
assign coef[29] = 17'b10000000011100110;
assign coef[30] = 17'b10000000111010110;
assign coef[31] = 17'b10000000101010111;
assign coef[32] = 17'b10000000000101111;
assign coef[33] = 17'b00000000011000000;
assign coef[34] = 17'b00000000011110110;
assign coef[35] = 17'b00000000010000010;
assign coef[36] = 17'b10000000000100111;
assign coef[37] = 17'b10000000010010000;
assign coef[38] = 17'b10000000010000110;
assign coef[39] = 17'b10000000000101000;
assign coef[40] = 17'b00000000000111100;
assign coef[41] = 17'b00000000001100111;
assign coef[42] = 17'b00000000001001001;
assign coef[43] = 17'b00000000000000001;
assign coef[44] = 17'b10000000001000100;
assign coef[45] = 17'b10000000001100110;
assign coef[46] = 17'b10000000001100000;
assign coef[47] = 17'b10000000001000011;
assign coef[48] = 17'b10000000000100011;
assign coef[49] = 17'b10000000000001101;
assign coef[50] = 17'b10000000000000010;
*/




// Коэффициенты КИХ-фильтра	часть процесса прямой код   8k 69 полоса ДЛЯ СИН_10 (синус с увеличивающейся частотой) !!!!!!!!!!
/*
assign coef[0] = 17'b10000000100001001;
assign coef[1] = 17'b10000000000010111;
assign coef[2] = 17'b10000000000100011;
assign coef[3] = 17'b10000000000110100;
assign coef[4] = 17'b10000000001000110;
assign coef[5] = 17'b10000000001010101;
assign coef[6] = 17'b10000000001011110;
assign coef[7] = 17'b10000000001011100;
assign coef[8] = 17'b10000000001001110;
assign coef[9] = 17'b10000000000110100;
assign coef[10] = 17'b10000000000001111;
assign coef[11] = 17'b00000000000100000;
assign coef[12] = 17'b00000000001010011;
assign coef[13] = 17'b00000000010001000;
assign coef[14] = 17'b00000000010111010;
assign coef[15] = 17'b00000000011100110;
assign coef[16] = 17'b00000000100001010;
assign coef[17] = 17'b00000000100100010;
assign coef[18] = 17'b00000000100101111;
assign coef[19] = 17'b00000000100101111;
assign coef[20] = 17'b00000000100100010;
assign coef[21] = 17'b00000000100001010;
assign coef[22] = 17'b00000000011100111;
assign coef[23] = 17'b00000000010111010;
assign coef[24] = 17'b00000000010000011;
assign coef[25] = 17'b00000000001000110;
assign coef[26] = 17'b00000000000000100;
assign coef[27] = 17'b10000000001000010;
assign coef[28] = 17'b10000000010000111;
assign coef[29] = 17'b10000000011001010;
assign coef[30] = 17'b10000000100000110;
assign coef[31] = 17'b10000000100111001;
assign coef[32] = 17'b10000000101011111;
assign coef[33] = 17'b10000000101111000;
assign coef[34] = 17'b00001111010000000;
assign coef[35] = 17'b10000000101111000;
assign coef[36] = 17'b10000000101011111;
assign coef[37] = 17'b10000000100111001;
assign coef[38] = 17'b10000000100000110;
assign coef[39] = 17'b10000000011001010;
assign coef[40] = 17'b10000000010000111;
assign coef[41] = 17'b10000000001000010;
assign coef[42] = 17'b00000000000000100;
assign coef[43] = 17'b00000000001000110;
assign coef[44] = 17'b00000000010000011;
assign coef[45] = 17'b00000000010111010;
assign coef[46] = 17'b00000000011100111;
assign coef[47] = 17'b00000000100001010;
assign coef[48] = 17'b00000000100100010;
assign coef[49] = 17'b00000000100101111;
assign coef[50] = 17'b00000000100101111;
assign coef[51] = 17'b00000000100100010;
assign coef[52] = 17'b00000000100001010;
assign coef[53] = 17'b00000000011100110;
assign coef[54] = 17'b00000000010111010;
assign coef[55] = 17'b00000000010001000;
assign coef[56] = 17'b00000000001010011;
assign coef[57] = 17'b00000000000100000;
assign coef[58] = 17'b10000000000001111;
assign coef[59] = 17'b10000000000110100;
assign coef[60] = 17'b10000000001001110;
assign coef[61] = 17'b10000000001011100;
assign coef[62] = 17'b10000000001011110;
assign coef[63] = 17'b10000000001010101;
assign coef[64] = 17'b10000000001000110;
assign coef[65] = 17'b10000000000110100;
assign coef[66] = 17'b10000000000100011;
assign coef[67] = 17'b10000000000010111;
assign coef[68] = 17'b10000000100001001;
*/











// Коэффициенты КИХ-фильтра	часть процесса прямой код   8k 41 ФВЧ
/*
assign coef[0] = 17'b00000000000010010;
assign coef[1] = 17'b00000000010110001;
assign coef[2] = 17'b10000000001101000;
assign coef[3] = 17'b10000000001100000;
assign coef[4] = 17'b10000000001010000;
assign coef[5] = 17'b10000000000001000;
assign coef[6] = 17'b00000000001011001;
assign coef[7] = 17'b00000000010010010;
assign coef[8] = 17'b00000000001101011;
assign coef[9] = 17'b10000000000011011;
assign coef[10] = 17'b10000000010110100;
assign coef[11] = 17'b10000000011110000;
assign coef[12] = 17'b10000000010000010;
assign coef[13] = 17'b00000000001111101;
assign coef[14] = 17'b00000000101111110;
assign coef[15] = 17'b00000000110110110;
assign coef[16] = 17'b00000000010010010;
assign coef[17] = 17'b10000000111101011;
assign coef[18] = 17'b10000010100000101;
assign coef[19] = 17'b10000011110011000;
assign coef[20] = 17'b00001011101101001;
assign coef[21] = 17'b10000011110011000;
assign coef[22] = 17'b10000010100000101;
assign coef[23] = 17'b10000000111101011;
assign coef[24] = 17'b00000000010010010;
assign coef[25] = 17'b00000000110110110;
assign coef[26] = 17'b00000000101111110;
assign coef[27] = 17'b00000000001111101;
assign coef[28] = 17'b10000000010000010;
assign coef[29] = 17'b10000000011110000;
assign coef[30] = 17'b10000000010110100;
assign coef[31] = 17'b10000000000011011;
assign coef[32] = 17'b00000000001101011;
assign coef[33] = 17'b00000000010010010;
assign coef[34] = 17'b00000000001011001;
assign coef[35] = 17'b10000000000001000;
assign coef[36] = 17'b10000000001010000;
assign coef[37] = 17'b10000000001100000;
assign coef[38] = 17'b10000000001101000;
assign coef[39] = 17'b00000000010110001;
assign coef[40] = 17'b00000000000010010;
*/



// Коэффициенты КИХ-фильтра	часть процесса прямой код   16k 39 ФВЧ
/*
assign coef[0] = 17'b10000000000110111;
assign coef[1] = 17'b00000000011000010;
assign coef[2] = 17'b00000000000011101;
assign coef[3] = 17'b10000000000010010;
assign coef[4] = 17'b10000000000100100;
assign coef[5] = 17'b10000000000101101;
assign coef[6] = 17'b10000000000110001;
assign coef[7] = 17'b10000000000110000;
assign coef[8] = 17'b10000000000101000;
assign coef[9] = 17'b10000000000011001;
assign coef[10] = 17'b10000000000000100;
assign coef[11] = 17'b00000000000010100;
assign coef[12] = 17'b00000000000101100;
assign coef[13] = 17'b00000000000111111;
assign coef[14] = 17'b00000000001001001;
assign coef[15] = 17'b00000000001000110;
assign coef[16] = 17'b00000000000110101;
assign coef[17] = 17'b00000000000011000;
assign coef[18] = 17'b10000000000001101;
assign coef[19] = 17'b10000000000110110;
assign coef[20] = 17'b10000000001011010;
assign coef[21] = 17'b10000000001110010;
assign coef[22] = 17'b10000000001111000;
assign coef[23] = 17'b10000000001101000;
assign coef[24] = 17'b10000000001000001;
assign coef[25] = 17'b10000000000000111;
assign coef[26] = 17'b00000000000111111;
assign coef[27] = 17'b00000000010000101;
assign coef[28] = 17'b00000000010111111;
assign coef[29] = 17'b00000000011011111;
assign coef[30] = 17'b00000000011011011;
assign coef[31] = 17'b00000000010101010;
assign coef[32] = 17'b00000000001001001;
assign coef[33] = 17'b10000000001000101;
assign coef[34] = 17'b10000000011110101;
assign coef[35] = 17'b10000000110111011;
assign coef[36] = 17'b10000001010000011;
assign coef[37] = 17'b10000001100111001;
assign coef[38] = 17'b10000001111001100;
assign coef[39] = 17'b10000010000101011;
assign coef[40] = 17'b00001101110110100;
assign coef[41] = 17'b10000010000101011;
assign coef[42] = 17'b10000001111001100;
assign coef[43] = 17'b10000001100111001;
assign coef[44] = 17'b10000001010000011;
assign coef[45] = 17'b10000000110111011;
assign coef[46] = 17'b10000000011110101;
assign coef[47] = 17'b10000000001000101;
assign coef[48] = 17'b00000000001001001;
assign coef[49] = 17'b00000000010101010;
assign coef[50] = 17'b00000000011011011;
assign coef[51] = 17'b00000000011011111;
assign coef[52] = 17'b00000000010111111;
assign coef[53] = 17'b00000000010000101;
assign coef[54] = 17'b00000000000111111;
assign coef[55] = 17'b10000000000000111;
assign coef[56] = 17'b10000000001000001;
assign coef[57] = 17'b10000000001101000;
assign coef[58] = 17'b10000000001111000;
assign coef[59] = 17'b10000000001110010;
assign coef[60] = 17'b10000000001011010;
assign coef[61] = 17'b10000000000110110;
assign coef[62] = 17'b10000000000001101;
assign coef[63] = 17'b00000000000011000;
assign coef[64] = 17'b00000000000110101;
assign coef[65] = 17'b00000000001000110;
assign coef[66] = 17'b00000000001001001;
assign coef[67] = 17'b00000000000111111;
assign coef[68] = 17'b00000000000101100;
assign coef[69] = 17'b00000000000010100;
assign coef[70] = 17'b10000000000000100;
assign coef[71] = 17'b10000000000011001;
assign coef[72] = 17'b10000000000101000;
assign coef[73] = 17'b10000000000110000;
assign coef[74] = 17'b10000000000110001;
assign coef[75] = 17'b10000000000101101;
assign coef[76] = 17'b10000000000100100;
assign coef[77] = 17'b10000000000010010;
assign coef[78] = 17'b00000000000011101;
assign coef[79] = 17'b00000000011000010;
assign coef[80] = 17'b10000000000110111;
*/

// Коэффициенты КИХ-фильтра	часть процесса прямой код   2k 15 ФВЧ
/*
assign coef[0] = 17'b10000000010011010;
assign coef[1] = 17'b00000000011011010;
assign coef[2] = 17'b10000000101010011;
assign coef[3] = 17'b00000000111011000;
assign coef[4] = 17'b10000001001011001;
assign coef[5] = 17'b00000001011000101;
assign coef[6] = 17'b10000001100001101;
assign coef[7] = 17'b00000001100100111;
assign coef[8] = 17'b10000001100001101;
assign coef[9] = 17'b00000001011000101;
assign coef[10] = 17'b10000001001011001;
assign coef[11] = 17'b00000000111011000;
assign coef[12] = 17'b10000000101010011;
assign coef[13] = 17'b00000000011011010;
assign coef[14] = 17'b10000000010011010;
*/


// Коэффициенты КИХ-фильтра	часть процесса прямой код   8k 115 полосовой
//*
assign coef[0] = 17'b10000000000010000;
assign coef[1] = 17'b10000000000000010;
assign coef[2] = 17'b10000000000111001;
assign coef[3] = 17'b00000000000000001;
assign coef[4] = 17'b00000000001010110;
assign coef[5] = 17'b00000000001110100;
assign coef[6] = 17'b00000000000111000;
assign coef[7] = 17'b10000000000100101;
assign coef[8] = 17'b10000000001000100;
assign coef[9] = 17'b10000000000011100;
assign coef[10] = 17'b00000000000000010;
assign coef[11] = 17'b10000000000011110;
assign coef[12] = 17'b10000000001000100;
assign coef[13] = 17'b10000000000100110;
assign coef[14] = 17'b00000000000100001;
assign coef[15] = 17'b00000000000111000;
assign coef[16] = 17'b00000000000010000;
assign coef[17] = 17'b00000000000000000;
assign coef[18] = 17'b00000000000110010;
assign coef[19] = 17'b00000000001011011;
assign coef[20] = 17'b00000000000101100;
assign coef[21] = 17'b10000000000101010;
assign coef[22] = 17'b10000000000111011;
assign coef[23] = 17'b10000000000001000;
assign coef[24] = 17'b10000000000000010;
assign coef[25] = 17'b10000000001001111;
assign coef[26] = 17'b10000000001111111;
assign coef[27] = 17'b10000000000110110;
assign coef[28] = 17'b00000000000111010;
assign coef[29] = 17'b00000000001000010;
assign coef[30] = 17'b10000000000000011;
assign coef[31] = 17'b00000000000000110;
assign coef[32] = 17'b00000000001111011;
assign coef[33] = 17'b00000000010110100;
assign coef[34] = 17'b00000000001000011;
assign coef[35] = 17'b10000000001010000;
assign coef[36] = 17'b10000000001001001;
assign coef[37] = 17'b00000000000010110;
assign coef[38] = 17'b10000000000010001;
assign coef[39] = 17'b10000000011001001;
assign coef[40] = 17'b10000000100001110;
assign coef[41] = 17'b10000000001010111;
assign coef[42] = 17'b00000000001110100;
assign coef[43] = 17'b00000000001001110;
assign coef[44] = 17'b10000000000111111;
assign coef[45] = 17'b00000000000101011;
assign coef[46] = 17'b00000000101110011;
assign coef[47] = 17'b00000000111010111;
assign coef[48] = 17'b00000000010000101;
assign coef[49] = 17'b10000000011001110;
assign coef[50] = 17'b10000000001010010;
assign coef[51] = 17'b00000000011000010;
assign coef[52] = 17'b10000000010010100;
assign coef[53] = 17'b10000010001010110;
assign coef[54] = 17'b10000011000001111;
assign coef[55] = 17'b10000000111100111;
assign coef[56] = 17'b00000010110100110;
assign coef[57] = 17'b00000100101110111;
assign coef[58] = 17'b00000010110100110;
assign coef[59] = 17'b10000000111100111;
assign coef[60] = 17'b10000011000001111;
assign coef[61] = 17'b10000010001010110;
assign coef[62] = 17'b10000000010010100;
assign coef[63] = 17'b00000000011000010;
assign coef[64] = 17'b10000000001010010;
assign coef[65] = 17'b10000000011001110;
assign coef[66] = 17'b00000000010000101;
assign coef[67] = 17'b00000000111010111;
assign coef[68] = 17'b00000000101110011;
assign coef[69] = 17'b00000000000101011;
assign coef[70] = 17'b10000000000111111;
assign coef[71] = 17'b00000000001001110;
assign coef[72] = 17'b00000000001110100;
assign coef[73] = 17'b10000000001010111;
assign coef[74] = 17'b10000000100001110;
assign coef[75] = 17'b10000000011001001;
assign coef[76] = 17'b10000000000010001;
assign coef[77] = 17'b00000000000010110;
assign coef[78] = 17'b10000000001001001;
assign coef[79] = 17'b10000000001010000;
assign coef[80] = 17'b00000000001000011;
assign coef[81] = 17'b00000000010110100;
assign coef[82] = 17'b00000000001111011;
assign coef[83] = 17'b00000000000000110;
assign coef[84] = 17'b10000000000000011;
assign coef[85] = 17'b00000000001000010;
assign coef[86] = 17'b00000000000111010;
assign coef[87] = 17'b10000000000110110;
assign coef[88] = 17'b10000000001111111;
assign coef[89] = 17'b10000000001001111;
assign coef[90] = 17'b10000000000000010;
assign coef[91] = 17'b10000000000001000;
assign coef[92] = 17'b10000000000111011;
assign coef[93] = 17'b10000000000101010;
assign coef[94] = 17'b00000000000101100;
assign coef[95] = 17'b00000000001011011;
assign coef[96] = 17'b00000000000110010;
assign coef[97] = 17'b00000000000000000;
assign coef[98] = 17'b00000000000010000;
assign coef[99] = 17'b00000000000111000;
assign coef[100] = 17'b00000000000100001;
assign coef[101] = 17'b10000000000100110;
assign coef[102] = 17'b10000000001000100;
assign coef[103] = 17'b10000000000011110;
assign coef[104] = 17'b00000000000000010;
assign coef[105] = 17'b10000000000011100;
assign coef[106] = 17'b10000000001000100;
assign coef[107] = 17'b10000000000100101;
assign coef[108] = 17'b00000000000111000;
assign coef[109] = 17'b00000000001110100;
assign coef[110] = 17'b00000000001010110;
assign coef[111] = 17'b00000000000000001;
assign coef[112] = 17'b10000000000111001;
assign coef[113] = 17'b10000000000000010;
assign coef[114] = 17'b10000000000010000;
//*/


// Коэффициенты КИХ-фильтра	часть процесса прямой код   8k 135 режекторный
/*
assign coef[0] = 17'b10000000001001101;
assign coef[1] = 17'b00000000010010101;
assign coef[2] = 17'b10000000000100011;
assign coef[3] = 17'b10000000000000111;
assign coef[4] = 17'b00000000000111010;
assign coef[5] = 17'b00000000000110111;
assign coef[6] = 17'b00000000000001000;
assign coef[7] = 17'b10000000000001100;
assign coef[8] = 17'b00000000000001011;
assign coef[9] = 17'b00000000000010111;
assign coef[10] = 17'b10000000000001000;
assign coef[11] = 17'b10000000000101110;
assign coef[12] = 17'b10000000000101000;
assign coef[13] = 17'b10000000000000011;
assign coef[14] = 17'b00000000000000111;
assign coef[15] = 17'b10000000000010011;
assign coef[16] = 17'b10000000000011010;
assign coef[17] = 17'b00000000000010001;
assign coef[18] = 17'b00000000000111100;
assign coef[19] = 17'b00000000000101110;
assign coef[20] = 17'b00000000000000011;
assign coef[21] = 17'b00000000000000001;
assign coef[22] = 17'b00000000000100110;
assign coef[23] = 17'b00000000000100101;
assign coef[24] = 17'b10000000000011011;
assign coef[25] = 17'b10000000001001101;
assign coef[26] = 17'b10000000000110010;
assign coef[27] = 17'b10000000000000001;
assign coef[28] = 17'b10000000000010000;
assign coef[29] = 17'b10000000001000011;
assign coef[30] = 17'b10000000000110010;
assign coef[31] = 17'b00000000000101010;
assign coef[32] = 17'b00000000001011111;
assign coef[33] = 17'b00000000000110001;
assign coef[34] = 17'b10000000000000001;
assign coef[35] = 17'b00000000000101010;
assign coef[36] = 17'b00000000001101100;
assign coef[37] = 17'b00000000001000000;
assign coef[38] = 17'b10000000000111110;
assign coef[39] = 17'b10000000001101111;
assign coef[40] = 17'b10000000000101001;
assign coef[41] = 17'b00000000000000000;
assign coef[42] = 17'b10000000001010111;
assign coef[43] = 17'b10000000010101000;
assign coef[44] = 17'b10000000001010001;
assign coef[45] = 17'b00000000001011010;
assign coef[46] = 17'b00000000001111110;
assign coef[47] = 17'b00000000000010101;
assign coef[48] = 17'b00000000000000110;
assign coef[49] = 17'b00000000010100111;
assign coef[50] = 17'b00000000100001010;
assign coef[51] = 17'b00000000001101000;
assign coef[52] = 17'b10000000010000110;
assign coef[53] = 17'b10000000010001010;
assign coef[54] = 17'b00000000000010110;
assign coef[55] = 17'b10000000000011100;
assign coef[56] = 17'b10000000101010110;
assign coef[57] = 17'b10000000111011100;
assign coef[58] = 17'b10000000010011000;
assign coef[59] = 17'b00000000011100110;
assign coef[60] = 17'b00000000010010001;
assign coef[61] = 17'b10000000010011101;
assign coef[62] = 17'b00000000010000011;
assign coef[63] = 17'b00000010000111111;
assign coef[64] = 17'b00000011000011110;
assign coef[65] = 17'b00000000111111010;
assign coef[66] = 17'b10000010111000110;
assign coef[67] = 17'b00001011001000111;
assign coef[68] = 17'b10000010111000110;
assign coef[69] = 17'b00000000111111010;
assign coef[70] = 17'b00000011000011110;
assign coef[71] = 17'b00000010000111111;
assign coef[72] = 17'b00000000010000011;
assign coef[73] = 17'b10000000010011101;
assign coef[74] = 17'b00000000010010001;
assign coef[75] = 17'b00000000011100110;
assign coef[76] = 17'b10000000010011000;
assign coef[77] = 17'b10000000111011100;
assign coef[78] = 17'b10000000101010110;
assign coef[79] = 17'b10000000000011100;
assign coef[80] = 17'b00000000000010110;
assign coef[81] = 17'b10000000010001010;
assign coef[82] = 17'b10000000010000110;
assign coef[83] = 17'b00000000001101000;
assign coef[84] = 17'b00000000100001010;
assign coef[85] = 17'b00000000010100111;
assign coef[86] = 17'b00000000000000110;
assign coef[87] = 17'b00000000000010101;
assign coef[88] = 17'b00000000001111110;
assign coef[89] = 17'b00000000001011010;
assign coef[90] = 17'b10000000001010001;
assign coef[91] = 17'b10000000010101000;
assign coef[92] = 17'b10000000001010111;
assign coef[93] = 17'b00000000000000000;
assign coef[94] = 17'b10000000000101001;
assign coef[95] = 17'b10000000001101111;
assign coef[96] = 17'b10000000000111110;
assign coef[97] = 17'b00000000001000000;
assign coef[98] = 17'b00000000001101100;
assign coef[99] = 17'b00000000000101010;
assign coef[100] = 17'b10000000000000001;
assign coef[101] = 17'b00000000000110001;
assign coef[102] = 17'b00000000001011111;
assign coef[103] = 17'b00000000000101010;
assign coef[104] = 17'b10000000000110010;
assign coef[105] = 17'b10000000001000011;
assign coef[106] = 17'b10000000000010000;
assign coef[107] = 17'b10000000000000001;
assign coef[108] = 17'b10000000000110010;
assign coef[109] = 17'b10000000001001101;
assign coef[110] = 17'b10000000000011011;
assign coef[111] = 17'b00000000000100101;
assign coef[112] = 17'b00000000000100110;
assign coef[113] = 17'b00000000000000001;
assign coef[114] = 17'b00000000000000011;
assign coef[115] = 17'b00000000000101110;
assign coef[116] = 17'b00000000000111100;
assign coef[117] = 17'b00000000000010001;
assign coef[118] = 17'b10000000000011010;
assign coef[119] = 17'b10000000000010011;
assign coef[120] = 17'b00000000000000111;
assign coef[121] = 17'b10000000000000011;
assign coef[122] = 17'b10000000000101000;
assign coef[123] = 17'b10000000000101110;
assign coef[124] = 17'b10000000000001000;
assign coef[125] = 17'b00000000000010111;
assign coef[126] = 17'b00000000000001011;
assign coef[127] = 17'b10000000000001100;
assign coef[128] = 17'b00000000000001000;
assign coef[129] = 17'b00000000000110111;
assign coef[130] = 17'b00000000000111010;
assign coef[131] = 17'b10000000000000111;
assign coef[132] = 17'b10000000000100011;
assign coef[133] = 17'b00000000010010101;
assign coef[134] = 17'b10000000001001101;
*/


endmodule